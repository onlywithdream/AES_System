//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18C
//Created Time: Fri Nov  4 20:53:53 2022

module Gowin_Boot_SP_8x2K_3 (dout, clk, oce, ce, reset, wre, ad, din);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [10:0] ad;
input [7:0] din;

wire [23:0] sp_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 8;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h43420240A002407D0085DCD8D4D0CCC8C4C0DCD8D4D0CCC8C4C000C04002020C;
defparam sp_inst_0.INIT_RAM_01 = 256'h478C51678F798505A77785854167CACE000041C05F5E5D5C4B4A494857565554;
defparam sp_inst_0.INIT_RAM_02 = 256'h08030403080406040A05080551678E0041678087877885A75067104732478932;
defparam sp_inst_0.INIT_RAM_03 = 256'h50475047A88F678E07A08F678E07A88F6750475047A88F678E67004706020202;
defparam sp_inst_0.INIT_RAM_04 = 256'h478F0F97C7009707FE009787872DFE4167FEAA8F678E876885A7AC855167A700;
defparam sp_inst_0.INIT_RAM_05 = 256'h85C78741672685C787416700470A0204020A0308030C050A0551676647C7FE07;
defparam sp_inst_0.INIT_RAM_06 = 256'h678F0028854167C787A885A72E41674167264167858586971C670F83C741672E;
defparam sp_inst_0.INIT_RAM_07 = 256'h24FE5067F75167C7FE416785009727874167FE2E416741678785A7002985C741;
defparam sp_inst_0.INIT_RAM_08 = 256'h67854167FEA02400854167FEA807E7470F2C18D6B1A0855167A75067C6275167;
defparam sp_inst_0.INIT_RAM_09 = 256'h85430707FE4167FEFC47F5FDA2F3FEFE07476B272724FE434967854167FE361F;
defparam sp_inst_0.INIT_RAM_0A = 256'hA7FB2041672A4167858546A72045A7A0208785A70085A72A1D67430707FE4167;
defparam sp_inst_0.INIT_RAM_0B = 256'h074767272720FEFD2A4967FD41678785A70085A72A4967416785416785858647;
defparam sp_inst_0.INIT_RAM_0C = 256'h804400FE0FFEFEFE101161008327F7272426CE80440F432726CE805400FEFEFE;
defparam sp_inst_0.INIT_RAM_0D = 256'h27FD4327FE9727A0074714FDCB272A2C2ED6804400472726CE804400472726CE;
defparam sp_inst_0.INIT_RAM_0E = 256'h270727FD43FD07FECB2797270727FD43FD0727FEFCFCFC18716100FEFEFDFC07;
defparam sp_inst_0.INIT_RAM_0F = 256'h27FD07FEC3FD972707274727FD0727FEFCFCFC18716100F8FE072726FECF2797;
defparam sp_inst_0.INIT_RAM_10 = 256'h6100FE02FE0802FEFE10116185FEFE10116100F8FE072726FEC3FD972707274B;
defparam sp_inst_0.INIT_RAM_11 = 256'hA0F707C707FE00FEFE87CE80540FFEFEFEFE43272ED68044FEC3274705FE1011;
defparam sp_inst_0.INIT_RAM_12 = 256'h26270DFC18716100FCFEFDFC07272EFDC3274327FDA026FDFCFC18716185F7FE;
defparam sp_inst_0.INIT_RAM_13 = 256'hCB4726270DFC18716100FCFEFEFE07278027C7FE87C727FE07272487A087C747;
defparam sp_inst_0.INIT_RAM_14 = 256'hFE0727804727FEFE000727807727FE0000FE0727804727FE0000FE072724C7FE;
defparam sp_inst_0.INIT_RAM_15 = 256'h0FFE0727804727FE0000FE0727804727FEFE000727000FFE0727804727FE0000;
defparam sp_inst_0.INIT_RAM_16 = 256'h0727804727FEFE000727807727FE0000FE0727804727FE0000FE072724C7FE00;
defparam sp_inst_0.INIT_RAM_17 = 256'h0439FEFE8785474327070DFC18D4716100807727FE0000FE072724C7FE000FFE;
defparam sp_inst_0.INIT_RAM_18 = 256'h8FFDFE0F8F47F7FE0F8F47478027F7FE0F8F47F7FE0F8F47470539FEFE878547;
defparam sp_inst_0.INIT_RAM_19 = 256'hFD0EFD000F8FFDFE0F8F47F7FE0F8F47478077072747F6FE0F8F47F7FEFE000F;
defparam sp_inst_0.INIT_RAM_1A = 256'hFD0F8F47C72704F787853E00072787853E00072704F787853E00072787853600;
defparam sp_inst_0.INIT_RAM_1B = 256'h270DFC18D6805450A08077072747C6FD000F8FFDFE0007278077072747C6FD00;
defparam sp_inst_0.INIT_RAM_1C = 256'hFEA024FEFEFDFC18716100FE8F00432726CE805400FEFEFDFC0727FD8547FE07;
defparam sp_inst_0.INIT_RAM_1D = 256'h0727FD4327FE9727FD04FDFDFC872C2ED4716100FCFEFEFE07278027C7216700;
defparam sp_inst_0.INIT_RAM_1E = 256'h4700FD0F8FC7206602FEFD00FD3F25FDE3672747FDFFFDA826476C27272CFDFC;
defparam sp_inst_0.INIT_RAM_1F = 256'hFCFC18D6805400F4FE07FDFC072726FEC32743FD400747FD35251502FEFD0047;
defparam sp_inst_0.INIT_RAM_20 = 256'h8EFD45FC0727F0252524FD07FDFC472726FEC39726FE9727FEA0260D272709FC;
defparam sp_inst_0.INIT_RAM_21 = 256'hFDFDFC872A2C2ED471615084FDFD91FD45F025FCFEFDFC0727F02525FD45F025;
defparam sp_inst_0.INIT_RAM_22 = 256'hFDFEFFFD45F025A824FEFBFDFEFE97270747DAFEFE072743FD0727FD0727FE02;
defparam sp_inst_0.INIT_RAM_23 = 256'h77331F1B17130F0B0703000000805400F02525F02583FD45E3272724FE3125F9;
defparam sp_inst_0.INIT_RAM_24 = 256'h7F85FBCF395BED84B3A01A75E29AC315F1CC26C0AFF07D762BC57B008008FFBB;
defparam sp_inst_0.INIT_RAM_25 = 256'hE994119EB90E668A1FC62E08EAA96D79625C0ADB1488DC733D17ECD221F58FA8;
defparam sp_inst_0.INIT_RAM_26 = 256'h050A008457DA5092CC16642549B2664E0B3D32CB448782FB9E38D5160F680DDF;
defparam sp_inst_0.INIT_RAM_27 = 256'h3CB04DEF9F0DA95F593133F4FE204B1B0E89716EE8852273CEEA416B03028F06;
defparam sp_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000028207D63267E61;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //Gowin_Boot_SP_8x2K_3
