//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18C
//Created Time: Fri Nov  4 20:52:42 2022

module Gowin_Boot_SP_8x2K_0 (dout, clk, oce, ce, reset, wre, ad, din);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [10:0] ad;
input [7:0] din;

wire [23:0] sp_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 8;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'hD2B20B00920B2AEF8BFEF6EEE6DED6CEC63E362E261E160E01068B00198B0B6F;
defparam sp_inst_0.INIT_RAM_01 = 256'hE70D830785EF104785EF07F103002201000100F6D6B696F6D6B696F2D2B292F2;
defparam sp_inst_0.INIT_RAM_02 = 256'h63136313631363136313631383E7850393E7C785AAEF4785A311638963E70963;
defparam sp_inst_0.INIT_RAM_03 = 256'h2385A385E70DE70085E709E70085E705A12385A385E709E705AD638963136313;
defparam sp_inst_0.INIT_RAM_04 = 256'hE78513F78503C7058323C785AA3E8383B1A3E709E785AAEF4785BDBE83478511;
defparam sp_inst_0.INIT_RAM_05 = 256'h07C78503713A07C785034D638963136313631363136313631383F7F4D785A3F4;
defparam sp_inst_0.INIT_RAM_06 = 256'h0785113A9C9347C7852587853A932103353E8361C7859C8A13F993D78583953A;
defparam sp_inst_0.INIT_RAM_07 = 256'h8583A3F7BA8307BA83137DBE8384C78583A9233A932103F5B58785793AF78503;
defparam sp_inst_0.INIT_RAM_08 = 256'hC78513BE8304908785933E83F491F4F4B4AA227901A9BE83478523E7843E83F4;
defparam sp_inst_0.INIT_RAM_09 = 256'hBEBAC705838305A3A3E7A103E7A103A3F4F78484F48583EF13C78513BE83EF13;
defparam sp_inst_0.INIT_RAM_0A = 256'h85AA3E83013E837D878587853E878504F5C5878585878536933EBAC7058383A9;
defparam sp_inst_0.INIT_RAM_0B = 256'h74F78404F4BA03833A933E8303F5918785E187853A93210361858339C785F487;
defparam sp_inst_0.INIT_RAM_0C = 256'h0501238313832323228272E7C4F784B4A40001053E93C4A4000145B2E78903A3;
defparam sp_inst_0.INIT_RAM_0D = 256'h988384212384C10029F7850344C4B4A400790501A3C4A40001050123C4A40001;
defparam sp_inst_0.INIT_RAM_0E = 256'h8AC4D883BA038983C498848AC4D883BA03C48D2323232322823201E383032384;
defparam sp_inst_0.INIT_RAM_0F = 256'hBA0389831803848AC498C4BA03C48D2323232322823201E30344F49183C49884;
defparam sp_inst_0.INIT_RAM_10 = 256'h729883338313B7232322827201232322823201E30344F491831803848AC498C4;
defparam sp_inst_0.INIT_RAM_11 = 256'hF7E1B7E186836383A30001453E9383E38323C4A40079053E83C4B4F4AE232282;
defparam sp_inst_0.INIT_RAM_12 = 256'hC4F4AE2322823201E383032384F49183C43D849883F4C1832323228272F78683;
defparam sp_inst_0.INIT_RAM_13 = 256'hB4F4C4F4AE2322823201E3830323C4E7C407BA8307C42523C4F447854785B4F4;
defparam sp_inst_0.INIT_RAM_14 = 256'h03C4E777C48D832383C4E7F7848583230303C4E757C4A583230303C4F407B583;
defparam sp_inst_0.INIT_RAM_15 = 256'h1303C4E7D7C4A583230303C4E757C485832383C47D231303C4E7F7C4AD832303;
defparam sp_inst_0.INIT_RAM_16 = 256'hC4E7A7C489832383C4E7F7848D83230303C4E777C4AD83230303C4F407BD8323;
defparam sp_inst_0.INIT_RAM_17 = 256'hAA3E8323E5C498C4C4F4AE2326068232E7F784B983230303C4F4079983231303;
defparam sp_inst_0.INIT_RAM_18 = 256'h85830393A4F7B9831394C4E7C4F7B98313E4F7B98313D484F4AA3E8323F1E4F4;
defparam sp_inst_0.INIT_RAM_19 = 256'h83638323138D830393E4F7B9831384C4E7F735C4B4F7B98313A4F7B983032313;
defparam sp_inst_0.INIT_RAM_1A = 256'h83138407C4F4F7A5A5AA3E83C4BE41AA3E83C4F4F7A545AA3E83C4BEE1AA3E83;
defparam sp_inst_0.INIT_RAM_1B = 256'hF4AE232279452201E7F735C494078D83231389830383C4E7F735C49407858323;
defparam sp_inst_0.INIT_RAM_1C = 256'h83F491832383232282721C03E213C4A4000145B201E3830323C44D03B42123C4;
defparam sp_inst_0.INIT_RAM_1D = 256'hC49883C40D23848A83638303A3B4A40006823201E3830323C4E7C407BA933E83;
defparam sp_inst_0.INIT_RAM_1E = 256'h1523831307B693FDB38383038384D503F7C47498830383F474F78484F4918323;
defparam sp_inst_0.INIT_RAM_1F = 256'h2323227945B201E3039D832384F48583843DB683B374988384F7913303836374;
defparam sp_inst_0.INIT_RAM_20 = 256'hEF03152344DF8444F4BA039983E3C4F4858318848A83C48A8304F784C4F4B623;
defparam sp_inst_0.INIT_RAM_21 = 256'h8303A3C4B4A40006822201EF0383EF031F8481E3830323449F8444B103DF8481;
defparam sp_inst_0.INIT_RAM_22 = 256'h0383EF039F8485F4C183EF038323449234E78D0323C498B683C43E03C4252363;
defparam sp_inst_0.INIT_RAM_23 = 256'h44001C1814100C08040003010045B24F84448F8485EF03E74484F4C1838485EF;
defparam sp_inst_0.INIT_RAM_24 = 256'h4543D04A6A205329521B09EB071804713436B79CADFACAFE30F2631B1001CC88;
defparam sp_inst_0.INIT_RAM_25 = 256'h9B69E1866148704BE81CBA656C8DE791C249E0DE46226064C45FCD10BC925150;
defparam sp_inst_0.INIT_RAM_26 = 256'hF78C90A75EFD6C5DD486726D76280842EEA654C4349B7C81BF3052B041BF8CCE;
defparam sp_inst_0.INIT_RAM_27 = 256'hC8AEA0932D196027B1881F789AC6FCAA6F1D471CE2E796F0974F3A01C1CAD0B8;
defparam sp_inst_0.INIT_RAM_28 = 256'h00000000000000000000000000000000000000000000000000000055E1BA1783;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //Gowin_Boot_SP_8x2K_0
