//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18C
//Created Time: Fri Nov  4 20:53:32 2022

module Gowin_Boot_SP_8x2K_2 (dout, clk, oce, ce, reset, wre, ad, din);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [10:0] ad;
input [7:0] din;

wire [23:0] sp_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 8;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h624200A28B0082E0000AFAF2EAE2DAD2CAC23A322A221A12068B01068B010000;
defparam sp_inst_0.INIT_RAM_01 = 256'h0D63E78523A03E9383E03A9347852606000B0B8B664626066646260662422202;
defparam sp_inst_0.INIT_RAM_02 = 256'hF700E700F700E700F700E700C7852307C78523933E003E830785E705F70963F7;
defparam sp_inst_0.INIT_RAM_03 = 256'hE709E715192385A3132D2385A3133D2385E709E705A92385A385E741F700E700;
defparam sp_inst_0.INIT_RAM_04 = 256'h83A3F7BA8307BA13F4E7A6933EB9F4478504E52385A33E803E83213AC7850301;
defparam sp_inst_0.INIT_RAM_05 = 256'hBE83938785A9BE83938785E741F700E700F700E700F700E700C785E30383F485;
defparam sp_inst_0.INIT_RAM_06 = 256'h8523017DBEC7850393393E83C1C78587858D878536933EBAC705F78D838785A1;
defparam sp_inst_0.INIT_RAM_07 = 256'h2384E78513F7850384C7853607BA8313478504F5C7858785AA3E8301D5BE8347;
defparam sp_inst_0.INIT_RAM_08 = 256'h8593C785F49123EF13C785F49DA3C983A3230006D1113AF785030785E383D785;
defparam sp_inst_0.INIT_RAM_09 = 256'h369C8A1374878504F4A163F481E3F4F48983E383032384F0C78593C785F4D087;
defparam sp_inst_0.INIT_RAM_0A = 256'h03F54D87851987853A932103DD81837523AA3E83013E835987859C8A13748785;
defparam sp_inst_0.INIT_RAM_0B = 256'h8583E383032304F4C1C785F48785AA3E83013E8385C78587853E87853A933E83;
defparam sp_inst_0.INIT_RAM_0C = 256'h8272E7C4F784B4A400010501A38313832323228272F79C832322822201E374F4;
defparam sp_inst_0.INIT_RAM_0D = 256'h83C49883F4BA031193E163449983232323228272E7058323228272E705832322;
defparam sp_inst_0.INIT_RAM_0E = 256'h038D83C498848AC49883BA038583C498848A8304C4B4A400794501F7C484F491;
defparam sp_inst_0.INIT_RAM_0F = 256'h03848AC498C4BA0385835803848A8304C4B4A400794501F7C48A8323C49883BA;
defparam sp_inst_0.INIT_RAM_10 = 256'h0501C4F78407FAB4A40001053EB4A400014501F7C48A8323C498C4BA038D8358;
defparam sp_inst_0.INIT_RAM_11 = 256'h3193E293E2F407F4F4AA228232F7C407C4F4DC8323228272B4D88303A3A40001;
defparam sp_inst_0.INIT_RAM_12 = 256'h2383A3A400794501F7C4C4F4918323C498839C83C42D23C4B4A40079053E93F4;
defparam sp_inst_0.INIT_RAM_13 = 256'hC5832383A3A400794501F744C4F48583238303843E8383F4C183239321938983;
defparam sp_inst_0.INIT_RAM_14 = 256'hC49D83230303C4F4078D83231303C4E717C49583230303C4E797C4B5832383C4;
defparam sp_inst_0.INIT_RAM_15 = 256'hF784B583230303C4E797C49583230303C4F4078583E7F784BD83230303C4E7B7;
defparam sp_inst_0.INIT_RAM_16 = 256'hA983230303C4F4078983231303C4E737C49D83230303C4E7B7C4BD832383C4E7;
defparam sp_inst_0.INIT_RAM_17 = 256'hA3E9D4F4AA3E83180393A3A40022794501231303C4E7E7C499832383C4E7F784;
defparam sp_inst_0.INIT_RAM_18 = 256'h35C4F4F7B98313E4F7B98303238313F4F7B9831394F7B98303A37DF4F4AA3E83;
defparam sp_inst_0.INIT_RAM_19 = 256'hC407B4E7F735C4B4F7B98313D4F7B98303231389830393F4F7B98313D4C4E7F7;
defparam sp_inst_0.INIT_RAM_1A = 256'hC4F7B9830383A393AA3EBD078D83AA3E590785832393AA3E5D078983AA3EF907;
defparam sp_inst_0.INIT_RAM_1B = 256'h83A3A400068292B21123138D830383C4E7F735C484078983231385830383C4E7;
defparam sp_inst_0.INIT_RAM_1C = 256'hC42D23C4F4C4A400790501C4D9879C832322822201F7C4C4F49183C4BE83F4C1;
defparam sp_inst_0.INIT_RAM_1D = 256'h9183849883F4BA0374F784C4F4B2232322794501F784C4F48583238303478507;
defparam sp_inst_0.INIT_RAM_1E = 256'h03E784F7B9838685F6C4740784110384A1B3038384C7844D2383E383032384F4;
defparam sp_inst_0.INIT_RAM_1F = 256'hB4A40006822201F7C48A74F4918323C498839C84F08A8384C10363F7C474E799;
defparam sp_inst_0.INIT_RAM_20 = 256'hFF8481F4C183EF038323449234E78D0323C498B683C43E03C42523638303A3C4;
defparam sp_inst_0.INIT_RAM_21 = 256'h84C4F4B6232323227945B23F8444FF8481EF03F78444F4C183EF03838481EF03;
defparam sp_inst_0.INIT_RAM_22 = 256'h84846F8485EF03152384EF8484F4BA039983E3C4F4858318848A83C48A8304F7;
defparam sp_inst_0.INIT_RAM_23 = 256'h66221E1A16120E0A0602000000822201EF0383EF03BF8485E3830323848D032F;
defparam sp_inst_0.INIT_RAM_24 = 256'h0233AA58BEB1002FD65A2CB280052331E5F79372A247C9AB676F77004004EEAA;
defparam sp_inst_0.INIT_RAM_25 = 256'h878E981D57F6B58B74B425AEF44E37E4AC243A0BB8904F197E4413F3DA38409F;
defparam sp_inst_0.INIT_RAM_26 = 256'h58D3AB9D46B948B65C98F6D1A224A1C3952394E943FF39D7A3A56ABB2D428928;
defparam sp_inst_0.INIT_RAM_27 = 256'hBBF53B9C7A4A7FEC10C7A85AC0793EBE62C51ADF373574E6CFDC118ABD0F1E45;
defparam sp_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000C14D60499;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //Gowin_Boot_SP_8x2K_2
