//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18C
//Created Time: Fri Nov  4 20:53:09 2022

module Gowin_Boot_SP_8x2K_1 (dout, clk, oce, ce, reset, wre, ad, din);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [10:0] ad;
input [7:0] din;

wire [23:0] sp_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 8;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'h4241A10240A08100C5DEDAD6D2CECAC6C2DEDAD6D2CECAC600C240007121A100;
defparam sp_inst_0.INIT_RAM_01 = 256'h2847C7506700064167002067A710CC110400005F5E5D5C4B4A49485756555443;
defparam sp_inst_0.INIT_RAM_02 = 256'h43078A074B078C0743078E07C75067C787004167870041678FAE82C740124746;
defparam sp_inst_0.INIT_RAM_03 = 256'h8F678E67504750F867504750F8675047A08F678E6750475047A08CC74B078D07;
defparam sp_inst_0.INIT_RAM_04 = 256'h5067F75167C7416747804167878544A7A00750475067870041672585C74167A0;
defparam sp_inst_0.INIT_RAM_05 = 256'h004167A7A085004167A7A08FC7470783074F07870747078E07C7FAFE516707FE;
defparam sp_inst_0.INIT_RAM_06 = 256'h5067A0854387004167264167858546A7A885A726416743070717F75167A6A885;
defparam sp_inst_0.INIT_RAM_07 = 256'h07278F0F97C7009727872185C7FE4167A6A024858546A7FB2C4167A8855167A7;
defparam sp_inst_0.INIT_RAM_08 = 256'h4967868647FE251D67858647FE47FDFCFC87D471002985C741678FFAFE87C7FE;
defparam sp_inst_0.INIT_RAM_09 = 256'h85971C6747A6A2030F004747F8474707FEFAFDFEFE0727008549678686470085;
defparam sp_inst_0.INIT_RAM_0A = 256'h678785A70085A72A1F674167854167FEFB2041672A4167858586971C6747A62A;
defparam sp_inst_0.INIT_RAM_0B = 256'hFEF4FDFEFE97274785858647A7FB284167204167858546A72845A72C4967FD41;
defparam sp_inst_0.INIT_RAM_0C = 256'h61008327F7272426CE804400FE0FFEFEFE10116185F7FEFE10116150EC474703;
defparam sp_inst_0.INIT_RAM_0D = 256'hC727FDA826FD4702A0004727FDFCFCFC1871610082FEFE1011610082FEFE1011;
defparam sp_inst_0.INIT_RAM_0E = 256'h07FECB2797270727FD43FD07FEC7279727FEA0262A2C2ED68054006127272CFD;
defparam sp_inst_0.INIT_RAM_0F = 256'h972707274B27FD07FEC3FD9727FEA0262A2C2ED68054004B27FDFE0727FD43FD;
defparam sp_inst_0.INIT_RAM_10 = 256'h44C327572787F72426CE8044002426CE8054004B27FDFE07274F27FD07FEC3FD;
defparam sp_inst_0.INIT_RAM_11 = 256'h0F8701870747DE070710116185F727C92726FDFC1871618547FEFEFE8726CE80;
defparam sp_inst_0.INIT_RAM_12 = 256'hFDFC872ED68054006827272CFDFC0727FD8FFD4327FE07272C2ED680440F0747;
defparam sp_inst_0.INIT_RAM_13 = 256'hFDFEFDFC872ED680540069272726FE00FE00972700FEA022FEFE21673167FDFE;
defparam sp_inst_0.INIT_RAM_14 = 256'h27FE0000FE072724C7FE000FFE0727804727FE0000FE0727804727FEFE000727;
defparam sp_inst_0.INIT_RAM_15 = 256'h7727FE0000FE0727804727FE0000FE072724C7FEA0807727FE0000FE07278047;
defparam sp_inst_0.INIT_RAM_16 = 256'hFE0000FE072724C7FE000FFE0727804727FE0000FE0727804727FEFE00072780;
defparam sp_inst_0.INIT_RAM_17 = 256'h8785470431FEC3FDFEFC872ED2D68054000FFE0727804727FEFE000727807727;
defparam sp_inst_0.INIT_RAM_18 = 256'h072747F6FE0F8F47F7FEFE00FD0F8F47F7FE0F8F47F7FEFEFE8785470531FEFE;
defparam sp_inst_0.INIT_RAM_19 = 256'h2784478077072747F6FE0F8F47F7FEFE000F8FFDFE0F8F47F7FE0F8F47478077;
defparam sp_inst_0.INIT_RAM_1A = 256'h27F7FE00FDFE0F8F3E8785C7FD843E8785C7FDFE0F8F3E8785C7FD84368785C7;
defparam sp_inst_0.INIT_RAM_1B = 256'hFC872ED471615400000F8FFDFE0007278077072747C6FD000F8FFDFE00072780;
defparam sp_inst_0.INIT_RAM_1C = 256'h27FE072726272ED68044C32707D7FEFE10116150006127272EFD3B25FDA826FD;
defparam sp_inst_0.INIT_RAM_1D = 256'hFDC327FDA024FD07470127270BFCFC18D680540068272726FE00FE00978787C7;
defparam sp_inst_0.INIT_RAM_1E = 256'hA08027F700978617C72647C727FD3D2502FEFDC327A727FEFDFCFEFDFC07272E;
defparam sp_inst_0.INIT_RAM_1F = 256'h2C2ED471615000422707472CFDFE0727FD8F972607FD4327FD0047672747FEFD;
defparam sp_inst_0.INIT_RAM_20 = 256'hF025A82AFD8AFDFDFE97270747DAFEFE072743FD0727FD0727FE02FDFDFC872A;
defparam sp_inst_0.INIT_RAM_21 = 256'h272709FCFCFC18D6805400F02525F0258BFD456327272AFD87FDFD3B2595FD45;
defparam sp_inst_0.INIT_RAM_22 = 256'h2525F02587FD45FE1727F0252524FD07FDFC472726FEC39726FE9727FEA0260D;
defparam sp_inst_0.INIT_RAM_23 = 256'h55111D1915110D0905010000006150F5FDFDFBFD45F025FCFDFEFE1727FD45F0;
defparam sp_inst_0.INIT_RAM_24 = 256'hF94DEF4CCBFCD1E33B6E83271296C7D8A53FFDA4D45982D7016B7C362002DD99;
defparam sp_inst_0.INIT_RAM_25 = 256'h1ED9F8C135033EBDDDA6787A56D5C895D306325EEE2A815DA7970CFFB69DA33C;
defparam sp_inst_0.INIT_RAM_26 = 256'hE4BCD88D15ED7065A468F88B5BD92EFA4CC27BDE8E2FE3F34036095499E6A155;
defparam sp_inst_0.INIT_RAM_27 = 256'hEB2AE0C9E5B551801207DDCDDBD25618B729F175F9ADACB4F2679113AF3F2CB3;
defparam sp_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000002169772B53;
defparam sp_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //Gowin_Boot_SP_8x2K_1
